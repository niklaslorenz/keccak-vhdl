library IEEE;
use IEEE.std_logic_1164.all;
use work.types.all;
use work.test_types.all;

package test_data is

end package test_data;